package fsm_pkg;

localparam a = 2'b00;
localparam b = 2'b01;
localparam c = 2'b10;
    
endpackage